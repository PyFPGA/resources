`define SECS 1
