entity Top0 is
end entity Top0;

entity Top1 is
end entity Top1;

-- entity Top2 is
-- end entity Top1;
