`define FREQ 10000000
