module Top0 ();
endmodule

module Top1 ();
endmodule

// module Top2 ();
// endmodule

/*
module Top3 ();
endmodule
*/
